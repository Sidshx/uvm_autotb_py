//File Name: uvm_test.sv
