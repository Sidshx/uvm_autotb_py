//File Name: fifo_sequence.sv
