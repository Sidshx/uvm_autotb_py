// Monitor: fifo_monitor.sv)
class fifo_monitor extends uvm_monitor;
    `uvm_object_utils(fifo_monitor)

endclass : fifo_monitor
