// Test: fifo_test.sv)
class fifo_test extends uvm_test;
    `uvm_object_utils(fifo_test)

endclass : fifo_test
