// Sequencer: fifo_seqr.sv
class fifo_sequencer extends uvm_sequencer#(fifo_seq_item);
    `uvm_object_utils(fifo_sequencer)

endclass : fifo_sequencer)
