//File Name: uvm_scoreboard.sv
