//File Name: uvm_sequencer.sv
