// Driver: fifo_driver.sv)
class fifo_driver extends uvm_driver#(fifo_seq_item);
    `uvm_object_utils(fifo_driver)

endclass : fifo_driver
