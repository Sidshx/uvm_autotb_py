// Sequence: fifo_seq.sv
class fifo_sequence extends uvm_sequence;
    `uvm_object_utils(fifo_sequence)

endclass : fifo_sequence)
