// Scoreboard: fifo_scoreboard.sv)
class fifo_scoreboard extends uvm_scoreboard;
    `uvm_component_utils(fifo_scoreboard)

endclass : fifo_agent
