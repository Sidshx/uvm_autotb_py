//File Name: fifo_sequencer.sv
