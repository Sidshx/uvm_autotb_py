//File Name: uvm_driver.sv
