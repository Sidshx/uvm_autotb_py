//File Name: uvm_sequence.sv
