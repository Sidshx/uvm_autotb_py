//File Name: fifo_tbench_top.sv
