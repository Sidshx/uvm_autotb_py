//File Name: uvm_env.sv
