// TBench Top: tbench_top.sv)
module tbench_top;
   
endmodule : tbench_top
