// Environment: fifo_env.sv)
class fifo_env extends uvm_env;
    `uvm_component_utils(fifo_env)

endclass : fifo_env
