//File Name: uvm_monitor.sv
