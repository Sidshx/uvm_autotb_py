//File Name: uvm_seq_item.sv
