//File Name: tbench_top.sv
