// TBench Top: uart_top.sv)
module tbench_top;
    import uvm_pkg::*;

    initial begin
        run_test();


    end

endmodule : tbench_top
