// Sequence Item: fifo_seq_item.sv
class fifo_seq_item extends uvm_sequence_item;
    `uvm_object_utils(fifo_seq_item)

endclass : fifo_seq_item) 
