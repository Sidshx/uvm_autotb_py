//File Name: uvm_agent.sv
