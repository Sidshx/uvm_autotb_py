// Agent: fifo_agent.sv)
class fifo_agent extends uvm_agent;
    `uvm_component_utils(fifo_agent)

endclass : fifo_agent
